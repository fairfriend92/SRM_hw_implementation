library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ***
-- this is a special counter: in case of overflow the counter is not reset,
-- instead it outputs the same number untill it receives a reset signal 
-- ***

entity counter is
  generic(width: integer);
  port(
    dataIn: in std_logic_vector (width-1 downto 0);
    clk, rst, dataEn: in std_logic;
    rco: out std_logic_vector (0 downto 0); -- rco stands for ripple carry out
                                            -- the type is vector to allow
                                            -- conversion from unsigned
    dout: out std_logic_vector (width-1 downto 0)
    );
end counter;

architecture behavioural of counter is
  signal rco_int: unsigned (0 downto 0):= "1"; 
  signal dout_int: unsigned (width-1 downto 0):= (others=> '0');
  -- these are internal signals used to do arithmetic
begin
  count: process(clk, rst)
  begin
    if(clk'event and clk= '1') then
      if(rst= '1') then -- if the chip is reset the output and the internal
        -- variables are zeroed out
        --report "counter: the counter has been reset";
        dout_int<= (others=> '0');
        rco_int<= "0";
      elsif(rst= '0') then
        if(rco_int= "0" and dataEn= '0') then -- if the data input is not
          -- enabled, counting reprises from the last number generated by the
          -- counter itself
          dout_int<= dout_int + 1;
          if(dout_int= 2**width - 2) then -- test the overflow condition and
            -- eventually raise the overflow flag
            rco_int<= "1"; 
          end if;
        elsif(rco_int= "1" and dataEN= '0') then
          dout_int<= dout_int; -- if the overflow flag has been raised counting
                               -- stops                                     
        elsif(dataEn= '1') then -- if the data input is enable counting starts
                                -- from the value of dataIn 
          --report "counter: dataIn has ben enabled";
          if(unsigned(dataIn)< 2**width-2) then -- if dataIn is exactly
            -- 2**width then we cannot count any further and the overflow
            -- condition has been met already
            dout_int<= unsigned(dataIn)+1;
            rco_int<= "0";
          else
            dout_int<= unsigned(dataIn);
            rco_int<= "1";
          end if;
        end if;
      end if;
    end if;
  end process count;
  dout<= std_logic_vector(dout_int);
  rco<= std_logic_vector(rco_int);
end architecture behavioural;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

-- ***
-- the following is a rudimentary lookup table (lut)
-- *** 

entity lut is
  generic(
    addr_width, data_width: integer;
    data_path: string -- among the generics we include the location of the file
                      -- used to initalize the rom
    );
  port(
    clk: in std_logic;
    addr: in std_logic_vector (addr_width-1 downto 0);
    data: out std_logic_vector (data_width-1 downto 0)
    );
end lut;

architecture behavioural of lut is

  subtype word is std_logic_vector (data_width-1 downto 0);
  type rom_type is array (integer range 0 to 2**addr_width-1) of word;
  file data_file: text is data_path;  -- this is the file used to initialize
                                      -- the rom
  signal rom: rom_type; 

begin
  -- in the following process we initialize the rom from a file. Since we can't
  -- read a file of std_logic_vectors firstly we read a file of ASCII
  -- characters, then we convert the strings in std_logic_vectors
  rom_init: process(clk)

  variable data_line: line;
  variable data_string: string (data_width-1 downto 0);
  variable i, j: integer;
  variable tmp: word; -- used to hold the vector while it's being translated
                      -- from a string before it's passed to the rom

  begin
    j:= 0;
    while not endfile(data_file) loop
      i:= 0;
      readline(data_file, data_line); -- here we read the line...
      read(data_line, data_string); -- ...and here we store it in a string
      while i< data_width loop -- in this loop we do the conversion for the i-th
                               -- character of the j-th string
        case data_string(i) is
          when '0'=> tmp(i):= '0';
          when '1'=> tmp(i):= '1';
          when others=> tmp(i):= '-';                          
        end case;
         i:= i+1;        
      end loop;
      --report "lut: j is " & integer'image(j);
      rom(j)<= tmp; -- we finally pass the vector to its rom location
      j:= j+1;
    end loop;

  end process rom_init;

  -- in the following process we serve the request of the stimulus
  -- according to the address provided

  addr_decod: process(clk)
  begin
    if(clk'event and clk= '1') then
      data<= rom(to_integer(unsigned(addr)));
    end if;
  end process addr_decod;

end architecture behavioural;

library ieee;
use ieee.std_logic_1164.all;

-- ***
-- in order to have a single lut for multiple synapses we need to access the
-- same lut multiple times in a single master clock period, therefore we need a
-- frequency divider
-- ***

library ieee;
use ieee.std_logic_1164.all;

entity freq_divider is
  generic(factor: integer);
  port(
    clk, rst: in std_logic;
    clk_div: out std_logic:= '0'
    );
end entity freq_divider;

architecture behavioural of freq_divider is
begin
  freq_division: process(clk, rst)

  variable index, counter: integer:= 0;

  begin
    if (clk'event and clk= '1') then
      if (rst= '1') then -- if the entity is reset the output and the internal
                         -- variables are zeroed out
        clk_div<= '0';
        index:= 0;
        counter:= 0;
      else
        if (index= factor) then -- after the appropriate number of clk periods
                                -- we assert the output
          clk_div<= '1';
          index:= 0;
          counter:= factor-1; -- this index counts the number of clk periods
                              -- that must elapse before clk_div goes down 
        else
          if (counter= 0) then -- if we have counted down to 0 it's time for
                               -- the clk_div to go down
            clk_div<= '0';
            index:= index+1;
          else
            clk_div<= '1'; -- keep clk_div high untill counter equals 0
            counter:= counter-1;
          end if;
         end if;
      end if;
    end if;
  end process freq_division;
end architecture behavioural;

-- ***
-- the next entity is a cluster of synapses. We group the synapses in order
-- to limit the number of luts and counters utilized. The number of synapses
-- we can group together is determined by the factor by which we divide the
-- frequency, therefore it is susceptible to physical limitations
-- ***

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.fixpt_lib.all;

entity clusterSyn is
  generic(numSyn, addrWidth: integer; dataPath_lut: string);
  -- the generics are:
  -- numSyn: number of synapses the cluster is made of.
  -- addrWidth: width of the address of each location of the lut
  -- dataPath_lut: path where the file used to initialize the lut is located
  port(
    clk, clk_div: in std_logic;
    spike: in std_logic_vector (numSyn-1 downto 0);
    current: out fixpt_word:= (scale=> 17, word=> (others=> '0'))
    );
  -- the ports are:
  -- clk, clk_div: divided and master clock, respectively
  -- spike: array of impulses, each representing a single spike.
  -- current: current response to the sum of the numSyn spikes
end entity;

architecture behavioural of clusterSyn is
  
  constant width: integer:= addrWidth;

  subtype addr is unsigned (width-1 downto 0);
  type addr_rom is array (numSyn-1 downto 0) of addr;

  component counter
    generic(width: integer);
    port(
      dataIn: in std_logic_vector (width-1 downto 0);
      clk, rst, dataEn: in std_logic;
      rco: out std_logic_vector (0 downto 0);
      dout: out std_logic_vector (width-1 downto 0)
      );
  end component counter;
  
  signal rst, dataEn: std_logic:= '0';
  -- signals with names such as "fanout_to_fanin" are striclty used to connect
  -- components through port mapping
  signal tmpAddr_to_dataIn: addr:= (others=> '0');
  signal dout_to_rom: std_logic_vector (width-1 downto 0):= (others=> '0');
 
  component lut 
    generic(
      addr_width, data_width: integer;
      data_path: string
      );
    port(
      clk: in std_logic;
      addr: in std_logic_vector (addr_width-1 downto 0);
      data: out std_logic_vector (data_width-1 downto 0)
      );
  end component lut;

  constant addr_width: integer:= width;
  constant data_width: integer:= 32; 
  constant data_path: string:= dataPath_lut;
  
  signal tmpAddr_to_lut: addr:= (others=> '0');
  signal lut_to_current: std_logic_vector(32-1 downto 0);

  signal spike_flag: std_logic:= '0';
  signal firstSpike_flag: std_logic_vector (numSyn-1 downto 0):= (others=> '0');
    
begin

-- in the following process the signal spike_flag is raised whenever the master
-- clock, that is clk_div, is high. This is done so that the  calculation of
-- the current response is carried out between subsequent clk_div periods. In
-- addition to that we also raise the flag firstSpike_flag when a spike is
-- detected for the first time. This will come in handy in the main process
  
  clockCheck: process(clk_div)
    variable index: integer:= 0;
  begin
    if(rising_edge(clk_div)) then
      spike_flag<= '1';
      while(index< numSyn) loop
        if(spike(index)= '1') then firstSpike_flag(index)<= '1'; end if;
        index:= index+1;
      end loop;
      index:= 0;
    elsif(falling_edge(clk_div)) then spike_flag<= '0'; end if;
  end process clockCheck;

  main: process(clk)

    variable index, flag, flag_2: integer:= 0;
    variable tmpAddr: addr_rom:= (others=> (others=> '0'));
    -- current_acc is an accumulator used to store temporarily the sum of the
    -- currents of each synapse
    variable current_acc: fixpt_word:= (scale=> 17, word=> (others=> '0'));
    variable lut_to_current_tmp: fixpt_word:=
      (scale=> 17, word=> (others=> '0'));
    variable lastAddress: std_logic_vector(addr_width-1 downto 0):=
      (others=> '1');

  begin

    -- every time the counter generates an address and every time a value for
    -- the current is read from the lut we have a delay of one clk period. The
    -- reason for this is that these two operations are carried out by two
    -- components, the aforementioned "counter" and "lut". 
    -- Therefore we cannot iterate the process over the synapses every new clk
    -- period but we have to wait for the delays to elapse. In order to do so
    -- we use the variable flag to internally count the clk periods  since the
    -- start of the computation. Essentialy we are defining a new clock period
    -- of length intermidiate between clk and clk_div.
    -- flag_2 is used to stop the computation if all the synapses have been
    -- served before falling_edge(clk_div)
    
    if(clk'event and clk= '1') then

      if(spike_flag= '1' and flag= 0 and flag_2= 0) then
        -- spike_flag tells us whether clk_div is high or low
        -- flag is used to count the number of clks elapsed since the rising
        -- edge of clk_div
        -- flag_2 signals the end of the computation
        flag_2:= 0;
        -- index is used to iterate over the synapses
        if(spike(index)= '1') then -- if the index-th synapse has received a
          -- spike the process of generating the addresses for the lut must
          -- start anew and therefore the counter must be reset
          rst<= '1';
        else
          -- otherwise the counting resumes from the last address, which has
          -- been previously stored in tmpAddr(index)
          rst<= '0';
          if(firstSpike_flag(index)= '1') then -- there is no need to abilitate
            -- counting process if the index-th synapse hasn't received a spike
            -- yet 
            dataEn<= '1';
            tmpAddr_to_dataIn<= tmpAddr(index);
          else dataEn<= '0'; end if;               
        end if;
        flag:= 1; -- this means: next time rising_edge(clk) is true, move to
                  -- the subsequent step of the computation     

      elsif(spike_flag= '1' and flag= 1 and flag_2= 0) then
        -- in this clk period we merely wait for the counter to generate an
        -- address
        flag:= 2; -- as before

      elsif(spike_flag= '1' and flag= 2 and flag_2= 0) then

        if(firstSpike_flag(index)= '1') then
          tmpAddr_to_lut<= unsigned(dout_to_rom); -- the address generated by
          -- the counter is passed to the lut
          tmpAddr(index):= unsigned(dout_to_rom); -- the address is also stored
          -- in this temporariry register to be fetched by the counter in case
          -- spike(index+1)= 0
        else
          tmpAddr_to_lut<= unsigned(lastAddress);
          tmpAddr(index):= unsigned(lastAddress);
        end if;
        flag:= 3; -- as before

      elsif(spike_flag= '1' and flag= 3 and flag_2= 0) then
        -- again in this clk period we're merely catchin up with the delay
        flag:= 4; -- as before

      elsif(spike_flag= '1' and flag= 4 and flag_2= 0) then

        -- if we have serverd all the synapses then we raise flag_2 and the
        -- computation doesn't go any further 
        if(index< numSyn-1) then index:= index+1; else flag_2:= 1; end if;

        -- the output of the lut is essentialy cast into a fixed point number
        lut_to_current_tmp.word:= signed(lut_to_current);

        -- the current of the index-th synapse is summed to those of the
        -- previous numSyn-(index-1) synapses
        current_acc:= sum_words(current_acc, lut_to_current_tmp);
        flag:= 0;

      elsif(spike_flag= '0' and flag= 0 and flag_2= 1) then        
        flag:= 1;
        -- finally the current is associated with the output
        index:= 0;
        current<= current_acc;
      elsif(spike_flag= '0' and flag= 1 and flag_2= 1) then
        current_acc.word:= (others=> '0');
        index:= 0;
        flag:= 0;
        flag_2:= 0;
      end if;

    end if;    
        
  end process main;

  counter_Syn: counter
    generic map(width=> width)
    port map(
      clk=> clk, dataEn=> dataEn, 
      dataIn=> std_logic_vector(tmpAddr_to_dataIn),
      dout=> dout_to_rom, rst=> rst
      );

  lut_Syn: lut
    generic map(
      addr_width=> addr_width, data_width=> data_width, data_path=> data_path
      )
    port map(
      clk=> clk, addr=> std_logic_vector(tmpAddr_to_lut),
      data=> lut_to_current
      );

end architecture behavioural;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.fixpt_lib.all;
use ieee.math_real.all;
use ieee.math_real.all;

entity transversalFilter is
  generic(order, dataWidth: integer; weightRom_path: string);
  port(
    clk, clk_div, enable: in std_logic;
    dataIn: in fixpt_word:= (scale=> 17, word=> (others=> '0'));
    dataOut: out fixpt_word:= (scale=> 17, word=> (others=> '0'))
    );
end entity transversalFilter;

architecture behavioural of transversalFilter is

  subtype data is signed (dataWidth-1 downto 0);
  type data_rom is array (order-1 downto 0) of data;

  file data_file: text is weightRom_path;
  signal weightRom: data_rom;
  signal spike_flag, first_clk_div: std_logic:= '0';

begin

  -- the weights of the filter are initialized from a txt file whose location
  -- can be passed through the generic weightRom_path
  
  rom_init: process(clk)

  variable data_line: line;
  variable data_string: string (dataWidth-1 downto 0);
  variable i, j: integer;
  variable tmp: data;
  
  begin
    j:= 0;
    while not endfile(data_file) loop
      i:= 0;
      readline(data_file, data_line); 
      read(data_line, data_string); 
      while i< dataWidth loop 
        case data_string(i) is
          when '0'=> tmp(i):= '0';
          when '1'=> tmp(i):= '1';
          when others=> tmp(i):= '-';                          
        end case;
         i:= i+1;        
      end loop;
      weightRom(j)<= tmp; 
      j:= j+1;
    end loop;
    
  end process rom_init;
  
  clockCheck: process(clk_div)    
  begin
    if(rising_edge(clk_div)) then spike_flag<= '1'; first_clk_div<= '1';
    elsif(falling_edge(clk_div)) then spike_flag<= '0'; end if;
  end process clockCheck;

  main: process(clk)

    variable index, index_2: integer:= 0;
    variable acc, weight_tmp, data_tmp, prod_tmp: fixpt_word:=
      (scale=> 17, word=> (others=> '0'));
    variable dataRom: data_rom:= (others=> (others=>'0'));
    variable dataIn_tmp: signed (dataWidth-1 downto 0);
    
  begin

    if(clk'event and clk= '1') then
      if(spike_flag= '1') then
        -- when the master clock is high we compute the sum of the products
        -- between the weights and the input
        index_2:= 0;
        while(index< order) loop -- the first order calculations must be handled
                                 -- separately
          weight_tmp.word:= weightRom(index); 
          if(index= 0) then
            dataIn_tmp:= dataIn.word; -- if order= 0 then the data is provided
                                      -- by the input
            acc:= prod_words(dataIn, weight_tmp); 
          else
            data_tmp.word:= dataRom(index-1); -- otherwise we take it from the
                                              -- past inputs store in dataRom
            prod_tmp:= prod_words(data_tmp, weight_tmp);
            acc:= sum_words(acc, prod_tmp);
          end if;
          index:= index+1;
        end loop;
      elsif(spike_flag= '0') then -- when the master clock is low we advance
                                  -- the input to the subsequent stage
        index:= 0;
        dataOut<= acc;
        while(index_2< order) loop
          if(index_2/= order-1) then 
            dataRom(order-1-index_2):= dataRom(order-1-index_2-1);
          else
            if(first_clk_div= '1' and enable= '1') then
              dataRom(0):= dataIn_tmp;
            elsif(first_clk_div= '1' and enable= '0') then
              -- if the transversal filter has not been enabled filtering halts
              -- and therefore no new value can be accepted
              dataRom(0):= (others=> '0');              
            else dataRom(0):= (others=> '0'); end if;                 
          end if;
          index_2:= index_2+1;
        end loop;
      end if;
    end if;

  end process main;
    
  end architecture behavioural;
    
        
                                                
                                                      
      
                                                      
                                                    
          
  
